typedef enum logic[2:0] {
    //TODO
}
packet_type
