//Including NoC
`include ../mesh_3x3/noc/toplevel.sv

//Including converters
`include ../converters/packet_collevtor.sv
`include ../converters/splitter.sv

